`ifndef FIFO_DEFINE_UVM
`define FIFO_DEFINE_UVM

`define DEPTH 16 //Depth of FIFO 
`define ADDR 4 //Address width 
`define WIDTH 8 //Data width 

`endif 

